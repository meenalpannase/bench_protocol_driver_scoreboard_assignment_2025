/************************************************************************
Author: Mirafra Technologies Pvt Limited
        By Meenal Pannase/Priya Ananthakrishnan
Filename:	Scoreborad.sv  
Date:   	29th Oct 2025
Version:	1.0
Description: Concept of scoreboard writing in UVM 
***************************************************************************/
//write scoreboard check for apb protocol, consider single master and single slave .

class scoreboard extends uvm_scoreboard
  //factory registration
  //declaration of ports from monitor/refrennce model
  //constructor
  //build phase
  //connect phase
  //run phase 
  //write scoreboard check here with expected and actual data
endclass
